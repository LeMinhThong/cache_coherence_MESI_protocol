`ifndef CACHE_UNITS_PKG_SV
`define CACHE_UNITS_PKG_SV

package cache_units_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  // agents
  `include "cache_vip_def.svh"
  `include "cache_type.svh"
  `include "cache_txn.svh"
  `include "cache_seqr.svh"
  `include "cache_drv_bfm.svh"
  `include "cache_drv.svh"
  `include "cache_mon.svh"
  `include "cache_agt.svh"

  // units
  `include "cache_model.svh"
  `include "cache_sb_base.svh"
  `include "cache_sb.svh"
  `include "cache_cov_def.svh"
  `include "cache_cov_cdreq.svh"
  `include "cache_cov_sureq.svh"
  `include "cache_cov.svh"
  `include "cache_env.svh"

  // Seqs
  `include "cache_base_seq.svh"
  `include "l1_req_seq.svh"
  `include "snp_req_seq.svh"

endpackage: cache_units_pkg

`endif
