`ifndef CACHE_VIP_DEF_SVH
`define CACHE_VIP_DEF_SVH

`define VIP_LINE_WIDTH      512   // 64 * 8
`define VIP_NUM_CACHE_LINE  1024
`define VIP_ADDR_WIDTH      64
`define VIP_DATA_WIDTH      32

`endif
