`ifndef CACHE_BASE_SEQ_SV
`define CACHE_BASE_SEQ_SV
`define THIS_CLASS cache_base_seq

class `THIS_CLASS extends uvm_sequence;
endclass: `THIS_CLASS

`undef THIS_CLASS
`endif
