`ifndef CACHE_TEST_PKG_SVH
`define CACHE_TEST_PKG_SVH

package cache_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh";

  `include "base_test.sv";
endpackage

`endif
