`ifndef CACHE_MEM_DEF_SVH
`define CACHE_MEM_DEF_SVH

`define LINE_WIDTH      64*8
`define NUM_CACHE_LINE  1024
`define ADDR_WIDTH      64
`define DATA_WIDTH      32

`endif
