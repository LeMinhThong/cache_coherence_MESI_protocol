`ifndef CACHE_MEM_IF_SV
`define CACHE_MEM_IF_SV


`endif
